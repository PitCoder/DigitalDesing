LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPARADOR IS
	PORT(A,B,C,D,SEL,REF: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 DISP1,DISP2: OUT STD_LOGIC_VECTOR(1 DOWNTO 0); 
		 DISP3: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPARADOR;

ARCHITECTURE ARQCOMPARADOR OF COMPARADOR IS
	BEGIN

	PROCESS(A, B, C, D, SEL, REF)
	VARIABLE TEMP1: STD_LOGIC_VECTOR(1 DOWNTO 0);
	VARIABLE TEMP2: STD_LOGIC_VECTOR(2 DOWNTO 0);
		BEGIN
				CASE SEL IS
					WHEN "00" => DISP1 <= A;
					WHEN "01" => DISP1 <= B;
					WHEN "10" => DISP1 <= C;
					WHEN OTHERS => DISP1 <= D;
				END CASE;
			
			TEMP1 := DISP1;

				IF REF=TEMP1 THEN
					TEMP2 := "100";
				ELSIF REF>TEMP1 THEN
					TEMP2 := "010";
				ELSE
					TEMP2 := "001";
			    END IF;

			DISP2 <= REF;

				IF TEMP2 = "100" THEN
					DISP3 <= "0101";
				ELSIF TEMP2 = "010" THEN
					DISP3 <= "1101";
				ELSE 
					DISP3 <= "0111";
				END IF;

	END PROCESS;			         
END ARQCOMPARADOR;